library ieee;
use ieee.std_logic_1164.all;
use work.eecs361_gates.all;
use work.eecs361.all;

entity datapath is
  port (
  );
end entity;

architecture structural of datapath is
begin
  
end architecture;
